module cpu (
	input clk, reset
);
	reg [31:0] rom [0:4095];

	always @(posedge clk) begin

	end
endmodule
